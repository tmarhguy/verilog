module tb_alu_comb;
    // TODO: Declare signals
    // TODO: Instantiate alu_comb
    // TODO: Create tasks for testing specific operations (exec_add, exec_sub)
    // TODO: Self-checking logic (assert output == expected)
endmodule
